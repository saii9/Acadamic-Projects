CIRCUIT C:\microwind2\Book on CMOS\invAmpli.MSK
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
Vin 11 0 PULSE(0.00 1.20 0.23N 0.02N 0.02N 0.23N 0.50N)
*
* List of nodes
* "inv3" corresponds to n�5
* "inv2" corresponds to n�7
* "inv1" corresponds to n�9
* "in" corresponds to n�11
*
* MOS devices
MN1 0 11 5 0 N1  W= 0.54U L= 0.12U
MN2 0 11 7 0 N1  W= 0.24U L= 0.12U
MN3 0 11 9 0 N1  W= 0.24U L= 0.12U
MP1 1 11 5 1 P1  W= 0.24U L= 0.12U
MP2 1 11 7 1 P1  W= 0.24U L= 0.12U
MP3 1 11 9 1 P1  W= 0.72U L= 0.12U
*
C2 1 0  1.358fF
C3 1 0  1.275fF
C4 1 0  1.275fF
C5 5 0  0.516fF
C7 7 0  0.437fF
C9 9 0  0.544fF
C11 11 0  1.122fF
*
*
* n-MOS BSIM4 :
* low leakage
.MODEL N1 NMOS LEVEL=14 VTO=0.40 U0=0.050 TOX= 3.5E-9 LINT=0.010U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.540 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  1.6 U0=0.050 UA=3.000e-15
+WINT=0.020U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.050
+XJ=0.150U NDEP=170.000e15 PCLM=1.100
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* p-MOS BSIM4:
* low leakage
.MODEL P1 PMOS LEVEL=14 VTO=-0.45 U0=0.018 TOX= 3.5E-9 LINT=0.010U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.540 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  1.6 U0=0.018 UA=3.000e-15
+WINT=0.020U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.050
+XJ=0.150U NDEP=170.000e15 PCLM=0.700
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* Transient analysis
*
.TEMP 27.0
.TRAN 0.30PS 2.00N
.PROBE
.END
